library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity test_vhdl is
	port(
		clk : in std_logic_vector(hi downto 0);
		rst : in std_logic
	);
end entity test_vhdl;

architecture RTL of test_vhdl is
	
begin

end architecture RTL;
