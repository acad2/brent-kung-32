library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity carry_generate_block is
	port(
		clk : in std_logic;
		rst : in std_logic
	);
end entity carry_generate_block;

architecture RTL of carry_generate_block is
	
begin

end architecture RTL;
