-----------------------------------------------------------------------------------------------------------------------
-- (C) Copyright 2012 <Company Name> All Rights Reserved
--
-- ENTITY:    entity_name
-- DEVICE:
-- PROJECT:
-- AUTHOR:    student
-- DATE:      2018 11:43:05 PM
--
-- ABSTRACT:  You can customize the file content form Templates "VHDL File"
--
-----------------------------------------------------------------------------------------------------------------------

entity entity_name is
	port(
		port_name : IN STD_LOGIC
	);
end entity entity_name;

architecture rtl of entity_name is
	--declarative part
begin
	--statement part
end architecture rtl;

-----------------------------------------------------------------------------------------------------------------------
--
-- REVISION HISTORY:
--
-----------------------------------------------------------------------------------------------------------------------
